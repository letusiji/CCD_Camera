module CCD_DEMO();
